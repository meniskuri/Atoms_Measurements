*
R22 N001 N007 0.005
R26 N008 N012 0.005
R30 N016 N015 0.005
R31 0 N003 1000000
C9 N013 N003 1e-009
L1 N002 N001 0.00015005
L2 N003 N002 1e-007
C17 N001 0 3e-010
C18 N002 0 2e-011
C19 N003 0 1e-010
C20 N002 N001 1.7e-009
C21 N003 N002 2e-012
R32 0 N013 0.001
R33 N002 N001 400
R34 N003 N002 100
L3 N010 0 2e-007
L11 N014 0 2e-007
L12 N005 N004 2e-007
L13 N006 N007 0.00011
L14 N011 N012 0.00011
L15 N018 N015 0.00011
C22 N007 N005 8e-008
C23 N012 N010 8e-008
C24 N015 N014 8e-008
R57 N012 N010 18
R58 N015 N014 18
R59 N007 N005 18
R60 N006 N005 0.01
R61 N011 N010 0.01
R62 N018 N014 0.01
L16 N009 N008 0.00015005
L17 N003 N009 1e-007
C25 N008 0 3e-010
C26 N009 0 2e-011
C27 N003 0 1e-010
C28 N009 N008 1.7e-009
C29 N003 N009 2e-012
R63 N009 N008 400
R64 N003 N009 100
L18 N017 N016 0.00015005
L19 N003 N017 1e-007
C30 N016 0 3e-010
C31 N017 0 2e-011
C32 N003 0 1e-010
C33 N017 N016 1.7e-009
C34 N003 N017 2e-012
R65 N017 N016 400
R66 N003 N017 100
V1 N004 0 AC 1 0 

.ac oct 64 40 50Meg 
.backanno 
.print I(V1) 

.end 
